.SUBCKT U2Tx%sy%s nWL nBL nIN
M1 n1 nIN 0 0 nmos W=500n L=50n
M2 n1 nWL nBL 0 nmosx%sy%s W=50n L=500n
.ENDS
